library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

entity logic is
	port (
		-------------------------------
		-- TODO
		-- Define Ports of logic entity
		-------------------------------
	);
end entity logic;

architecture behav of logic is

	-------------------------------
	-- TODO (if required)
	-- Define additional signals
	-------------------------------

begin

	-------------------------------
	-- TODO
	-- Define logic behavior
	-------------------------------

end behav;

