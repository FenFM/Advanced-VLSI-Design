library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


entity hazard_detection_unit is
    port(
        
    );
end hazard_detection_unit;


architecture behavior of hazard_detection_unit is


begin


end behavior;
